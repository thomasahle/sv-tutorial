module top;
  initial begin
    // TODO: $display("HELLO WORLD");
  end
endmodule
