module top;
  initial begin
    $display("HELLO WORLD");
  end
endmodule
